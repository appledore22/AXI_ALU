module axi_fifo(clk,reset,wdata,wvalid,wready,rvalid,rdata,rready);
  
  input clk;
  input reset;
  
  // write data channel
  input [7:0] wdata;
  input wvalid;
  output reg wready;	
  
  // read data channel
  output reg rvalid;
  output reg [7:0] rdata;
  input rready;
  
  reg full;
  reg empty;
  
  reg [7:0] mem [8];
  reg [2:0] wptr;
  reg [2:0] rptr;
  
  assign wready = ~full;	// fifo not full. So ready to take write data
  assign rvalid = ~empty;	// fifo not empty. So output data is valid until fifo not empty to send data
  
  always@(posedge clk)
    begin
      if(reset)
        begin
          wptr <= 0;
          rptr <= 7;
          full <= 0;
          empty <= 1;
        end
      else
        begin
            if(wvalid && wready)
              begin
                mem[wptr] <= wdata;
                empty <= 0;
                if(wptr == (rptr-1) || (wptr == 7 && rptr == 0))
                	wptr <= wptr;
                else
                  wptr <= wptr +1;
              end          	
          	if(wptr == (rptr-1) || (wptr == 7 && rptr == 0))
              begin
              	full <= 1;
                empty <= 0;
                
              end
          	if(rptr == wptr)
              begin
               empty <= 1;
               full  <= 0;
              end         	
        end      
    end 
  
  always@(negedge clk)
    begin
      if(!empty)
              begin
                rdata <= mem[rptr];
                if(rready)
                	rptr <= rptr + 1;
              end
          
    end
  
endmodule
